`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    18:01:56 04/27/2016 
// Design Name: 
// Module Name:    MUX_salida 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module MUX_salida(
    input [8:0] in_inicio,
    input [8:0] in_lectura,
    input [8:0] in_escritura,
    input Sel_in,
    input Sel_rd,
    input Sel_wr,
    inout [8:0] RTC
    );


endmodule
