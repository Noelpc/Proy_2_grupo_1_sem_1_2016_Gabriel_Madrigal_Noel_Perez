`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:46:12 04/19/2016 
// Design Name: 
// Module Name:    DecoDir_countDir 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DecoDir_countDir(
    );

Dir_escritura instance_name (
    .binary_in(binary_in), 
    .decoder_out(decoder_out), 
    .EN(EN)
    );



endmodule
